library verilog;
use verilog.vl_types.all;
entity ULA_JUAN_THALES_vlg_vec_tst is
end ULA_JUAN_THALES_vlg_vec_tst;
