LIBRARY	IEEE;
USE IEEE.std_logic_1164.all;

ENTITY seg7_2 IS
  PORT(
  entrada: in std_logic_vector(3 downto 0);
  s: out std_logic_vector(13 downto 0)
  );
END seg7_2;

ARCHITECTURE arq_seg7_2 OF seg7_2 IS
BEGIN 
  WITH entrada SELECT
  
  s <=	"11111111000000" WHEN "0000", -- 00
			"11111111111001" WHEN "0001", -- +1
			"11111110100100" WHEN "0010", -- +2
			"11111110110000" WHEN "0011", -- +3
			"11111110011001" WHEN "0100", -- +4
			"11111110010010" WHEN "0101", -- +5
			"11111110000010" WHEN "0110", -- +6
			"11111111111000" WHEN "0111", -- +7
			"01111110000000" WHEN "1000", -- -8
			"01111111111000" WHEN "1001", -- -7     
			"01111110000010" WHEN "1010", -- -6
			"01111110010010" WHEN "1011", -- -5
			"01111110011001" WHEN "1100", -- -4
			"01111110110000" WHEN "1101", -- -3
			"01111110100100" WHEN "1110", -- -2
			"01111111111001" WHEN "1111"; -- -1
end arq_seg7_2;